`include "config.vh"

module top
(
    input        clk,
    input        reset_n,
    
    input  [3:0] key_sw,
    output [3:0] led,

    output [7:0] abcdefgh,
    output [3:0] digit,

    output       buzzer,

    output       hsync,
    output       vsync,
    output [2:0] rgb
);

    wire reset = ~ reset_n;

    assign abcdefgh  = 8'hff;
    assign digit     = 4'hf;
    assign buzzer    = 1'b0;
    assign hsync     = 1'b1;
    assign vsync     = 1'b1;
    assign rgb       = 3'b0;

    // Exercise 1: Free running counter.
    // How do you change the speed of LED blinking?
    // Try different bit slices to display.

    /* reg [31:0] cnt;
    
    always @ (posedge clk or posedge reset)
      if (reset)
        cnt <= 32'b0;
      else
        cnt <= cnt + 32'b1;

    assign led = ~ cnt [30:27]; */

    // Exercise 2: Key-controlled counter.
    // Comment out the code above.
    // Uncomment and synthesize the code below.
    // Press the key to see the counter incrementing.
    //
    // Change the design, for example:
    //
    // 1. One key is used to increment, another to decrement.
    //
    // 2. Two counters controlled by different keys
    // displayed in different groups of LEDs.

    

    wire key = key_sw [0];
    reg key_r;
    always @ (posedge clk or posedge reset)
      if (reset)
        key_r <= 1'b0;
      else
        key_r <= key;
    wire key_pressed = ~ key & key_r;
	 
	 wire key2 = key_sw [3];
    reg key_d;
    always @ (posedge clk or posedge reset)
      if (reset)
        key_d <= 1'b0;
      else
        key_d <= key2;
    wire key_d_pressed = ~ key2 & key_d;

	 reg inc_dec;
	 always @ (posedge clk or posedge reset)
		if (reset)
			inc_dec <= 1'b0;
		else if (key_d_pressed)
			inc_dec <= inc_dec + 1'b1;
			
    reg [3:0] cnt;
    always @ (posedge clk or posedge reset)
      if (reset)
        cnt <= 4'b0;
      else if (key_pressed & ~ inc_dec)
        cnt <= cnt + 4'b1;
		else if (key_pressed & inc_dec)
			cnt <= cnt - 4'b1;

    assign led = ~ cnt;

    

endmodule
